{{ _header }}

    tran tr(PLUS, MINUS);

endmodule
